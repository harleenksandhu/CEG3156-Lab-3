library ieee;
use ieee.std_logic_1164.all;

entity pipeline_datapath is
	port(GClk, GReset: in std_logic);
	
end pipeline_datapath;


architecture rtl of pipeline_datapath is 



begin 


end rtl;